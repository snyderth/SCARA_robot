module	SinDeg(input	signed	[7:0]	data_in
			output real data_out);


		case(data_in):
			-90: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001100011000001011100011110000011000000110000010111000111100000110000001100000101110001111000001100000011000001011100011110000011000000110000010111000111100000110000001100000101110001111000001100000011000000100111;
			-89: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001011100011110000110011001100101010111000111100001100011001100000101110001111000001110010011011101011100011110000110011000110101010111000111100001100001011001100101110001111000001110000110000100100111;
			-88: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001011100011110000110011001100010010111000111100000110000001100100111100001011100011110000110001001100110010111000111100000110000001101010110011100100111;
			-87: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001011100011110000110011000110100010111000111100001100011001101010101110001111000011001010110010001011100011110000011000100110010010111000111100001100101001101100101110001111000001100010110010000100111;
			-86: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001011100011110000110010101100011010111000111100000110000011000100111000101110000010111000111100001100110011001100101110001111000011001100011011000100111;
			-85: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001011100011110000110010100110000010111000111100001100100001100110101110001111000011000100011010001011100011110000011000100111000010111000111100000110001001101010101110001111000011000010011001000100111;
			-84: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001011100011110000110010000110011010111000111100000110001011001100101110001111000001110010011010001011100011110000110011000111000011001110101110001111000011000110011011000100111;
			-83: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001011100011110000110001100110010010111000111100001100110001100000010010101011100011110000110000100110010001111100101110001111000001110000110001000100111;
			-82: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001011100011110000110001000110000010001100101110001111000011000010011100100110000010111000111100000111001001101000111100100100111;
			-81: data_out = 011000100010011101011100011110000110001001100110010111000111100001100101011001100101110001111000001110010110001000100100010111000111100000111001001101000010111101011100011110000110010100110100010111000101110000100111;
			-80: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001011100011110000011100000110011010111000111100000111000011000100101110001111000001110000110001101011100011110000011100000110001010111000111100000110001011000110101110001111000001100010011011100100111;
			-79: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001101001011111010110100100111000010111000111100001100010001101100101110001111000011000110011001000100111;
			-78: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001001100010111000111100001100110011000110011001001111010010111000111100000110000001100000101110001111000001101110110011000100111;
			-77: data_out = 011000100010011101011100011110000110001001100110010111000111100001100101011001100010111001011100011011100010000101001110010111000111100000111000001101110101110001111000001100000110011000100111;
			-76: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110011001011100011110000011000001100011010111000111100001100001001110010101110001111000001110010110011001111001010111000111100001100010011000010010010100100111;
			-75: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110010101011100011110000110010100111000010111000111100001100100011001000100011101001000010111000111100001100010011001100101110001111000001100010011010100100111;
			-74: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110010101011100011110000110001100110010010111000111100001100001001101110101110001111000011001010011001101011110011110110101110001111000001110000011000000100111;
			-73: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110010101011100011110000011100101100001010111000111100000110000011000110110111001111011010111000111100001100100011000100101110001111000001100010110011000100111;
			-72: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110010101101111010111000111100000110000011001010101110001111000001100010011001101000100010101000101110001111000011001100110011000100111;
			-71: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110010101000001010111000111100001100010001100000010101101011100011110000110011001100101010111000111100001100010001101000101110001111000011000110110000100100111;
			-70: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110010101011100011110000011000100110001010111000111100001100110001101100100001001010010001011010101110001111000001100010110001000100111;
			-69: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110010001011100011110000110010001100110010111000111100001100101001101000101110001111000001100000110010101011100011110000110011001100110010111000111100001100010001110000101110001111000001100000011010100100111;
			-68: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110010001011100011110000110000101100010011111010111100101011100011110000011100100110111010111000111100001100011011000100101100000100111;
			-67: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110010001110100010111000111100001100011001101100101110001111000001110010011100000101100011001100110111000100111;
			-66: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110010000111011010111000111100001100011001100110101110001111000011000010110010101011100011110000110011001100110010111000111100000110111011001100101110001111000001110010011010100100111;
			-65: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110010001011100011110000011000000110000011110010011000000101101010111000111100001100100001101110110011100100111;
			-64: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110001101011100011110000110001100110010010111000111100001100101011000100101110001111000011000100110001001010110001110000101110001111000011000110110000100100111;
			-63: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110001101011100011110000011100000110011001000000101110001111000001100010110010000111101001011000110110000100111;
			-62: data_out = 0110001000100010010111000111100001100010011001100101110001111000011001010110001101000001010111000111100000110001011000100100111101101101001001110101110001111000001100000011011100100010;
			-61: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110001001011100011110000110011001100011010111000111100001100101001100100111011101011100011110000110010000110011001110010101110001111000011000110011011000100111;
			-60: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110001001011100011110000110001000110110011110100101110001111000011001010011100001011000010011000101110001111000011000010110000100100111;
			-59: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110001001101101010111000111100001100101011000010101110001111000001100010110010101110110010111000111100001100101011000010101110001111000011001000110010000100111;
			-58: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110001000100011001101010101110001111000011000110011001001011100011110000110001101100100010111000111100001100001001110010100010100100111;
			-57: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110000101011100011110000110010000110110011000110101110001111000011000010011100001011100011110000110000101100101001011110101110001111000011001000110001000100111;
			-56: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110000101011100011110000011100000110111011110010101110001111000011000110110010001011100011110000110000100111000010111000111100001100101011001010101110001111000011000010011010100100111;
			-55: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010110000100110110011111100101100101011100011110000011000100110101010111000111100000111000001101110100011100100111;
			-54: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011100101011100011110000110010100110011011101110101110001111000001110010110001001011100011110000011100100110111010111000111100001100110001101000101110001111000011000010011100000100111;
			-53: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011100101011100011110000011100001100101011011000101110001111000001100000110010101011100011110000110000100110010011110100101110001111000001100010011010000100111;
			-52: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011100100110111011000100101001101011100011110000110011000110100011000110101110001111000011001000011001000100111;
			-51: data_out = 0110001000100010010111000111100001100010011001100101110001111000011001010011100001011100011110000110010001100101011000010011010101011100011110000011000100110101010111000111100001100001001100110010011100100010;
			-50: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011100001011100011110000011100000110011011011110101110001111000011000010011001001011100011110000110001101100110010100000011100100100111;
			-49: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011100000100110010111000111100000111001001101000101110001111000011000100011010001011100011110000110000100110001010111000111100000110001011000110011011100100111;
			-48: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011011101011100011110000110001100110111010111000111100001100100001101110101110001111000011000010011100000110011010111000111100001100010011001010101110001111000011000110011000100100111;
			-47: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011011101100111001111110101110001111000011001010011000001011100011110000110001100111000011010010101110001111000001110000011001000100111;
			-46: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011011101011100011110000011000000110100010111000111100001100100001101000101110001111000011001010011011001011100011110000110000100110101010011010011100000100111;
			-45: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011011001011100011110000110000100110000010111000111100000111001011001010110011001011100011110000011011101100110001110110101110001111000011000110110001100100111;
			-44: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011011000111010010111000111100001100001001101000011000001011100011110000110010100110000011100110101110001111000001100010011000000100111;
			-43: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011010101011100011110000110010000110010010111000111100001100101011001010011100101011100011110000011100001100011010111000111100000111001011000110010101100100111;
			-42: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011010101101001010111000111100000111000001101000101110001111000001110010011011001011100011110000110010100110010010111000111100000110000011000100101110001111000011001000011100000100111;
			-41: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011010001011100011110000110011001100101011011110101110001111000001110000011000100111000010011110101110001111000011001000011001100100111;
			-40: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011010001011100011110000011100100110001010111000111100001100010001101110101001000111100010111000111100000110001001101100101110001111000001100010110001100100111;
			-39: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011010000100011011001000101110001111000001110000011010001001000011110100101110001111000011000100110010000100111;
			-38: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011001101011100011110000110001000110011010111000111100000110111011001100101110001111000011000100011000101011100011110000110001001100100010111000111100001100011001110010011100000100111;
			-37: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011001101000010010111000111100000110001001100010101110001111000001110010011010001010101010111000111100001100010011001010101110001111000011000100011011000100111;
			-36: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011001001011100011110000110001101100110001000110101110001111000001100000011010001110101010110100101111000100111;
			-35: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011001001011010010111000111100001100010011000110101110001111000011001100011100001111100010010010111100000100111;
			-34: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011000101011100011110000110010100110100010111000111100001100101001110000101110001111000001110000011010001011100011110000011000100110001010111000111100001100110011001000101110001111000001100010011001100100111;
			-33: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011000101101101010111000111100001100001011001010101110001111000011001000011011101110000011101110101110001111000001100010110010000100111;
			-32: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011000001011100011110000110011000110101010111000111100000110001001110010011111001011100011110000110000101100011010111000111100001100100011001000010101000100111;
			-31: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001010011000001111011001100010010000001011100011110000110011001100100010111000111100001100100011001100101110001111000001100010011001100100111;
			-30: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000110011001011100011110000110011001100110010111000111100001100110011001100101110001111000011001100110011001011100011110000110011001100110010111000111100001100110011001100101110001111000011001100110011000100111;
			-29: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000110011001011100011110000011000000110111010111000111100000110001011001010101110001111000011001010110010001011100011110000110010101100110010111000111100001100001001100000101110001111000011001010110010000100111;
			-28: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000110010101011100011110000011000001100010010111000111100001100100001100100111010000100100010100000111100100100111;
			-27: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000110010001011100011110000011000001100101001011100010101101000100010111000111100001100100011001010101110001111000001100000011000000100111;
			-26: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000110001101011100011110000011000001100101010001010101110001111000011001000110000101011100011110000110001001100101010111000111100000110000001101010101110001111000011000110011100000100111;
			-25: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000110001001011100011110000011000001100011001011010111011100110111010111000111100000111001001110000101001100100111;
			-24: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000110000101011100011110000011000000110111010111000111100001100110001110010010000101011100011110000011000000110110010111000111100000110001011000010101110001111000011001000011000000100111;
			-23: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000011100101011100011110000011000000110001010111000111100001100010011001000010001001011100011110000011100100111000010111000111100001100110011001100101110001111000011000010110000100100111;
			-22: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000011011101011100011110000110011000111001010111000111100000111000011001000101110001111000011001010110010101011100011110000110010100110101010111000111100000111001001101100101110001111000001110000011000100100111;
			-21: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000011011001011100011110000110010101100110010111000111100000111000001100000101110001111000001100010110011001011100011110000110001101100101010111000111100001100100001100110011110000100111;
			-20: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000011010101011100011110000110010100110011010111000111100001100001001110000111010001011100011110000011100001100001010111000111100000110000011000100101110001111000011001100011010100100111;
			-19: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000011010001011100011110000110010000110110010111000111100000110001011000100101110001111000011001000011000001011100011110000011000000110000010111000111100001100011011001000101110001111000011001000110001000100111;
			-18: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000011001101011100011110000110001100110110010111000111100001100101011001100011011100101111010111000111100001100101001110010100111100100111;
			-17: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000011001001011100011110000110001000110110001101110101110001111000011000110110011001011100011110000011100000110011010111000111100001100100001101010101110001111000011000110011100000100111;
			-16: data_out = 011000100010011101011100011110000110001001100110010111000111100001100100001100010101110001111000011000010011010001011100011011100101110001111000011001000110010000110010010111000111100000111000011001010010100100100111;
			-15: data_out = 0110001000100111010111000111100001100010011001100101110001111000011001000011000001011100011110000011100100110000011111010101110001111000011000110011000101011100011110000011100100110011010111000111100000110000001101100101110001111000001110010011000000100111;
			-14: data_out = 0110001000100111010111000111100001100010011001100101110001111000011000110110010101011100011110000110011000110111010010110101110001111000011001100011001001011100011110000110010100110100010111000111100001100010001110010101110001111000001100010110010000100111;
			-13: data_out = 0110001000100111010111000111100001100010011001100101110001111000011000110110001101011100011110000110001101100010001100100011011001011100011110000110001101100100010111000111100001100011001101100111010100100111;
			-12: data_out = 0110001000100111010111000111100001100010011001100101110001111000011000110110000101011100011110000011100101100011010111000111100001100100001110010101110001111000011000010110001101000010010110000101110001111000011001100011010100100111;
			-11: data_out = 0110001000100111010111000111100001100010011001100101110001111000011000110011100001101100011011010101110001111000011001000110010001110110011000100100111100100111;
			-10: data_out = 0110001000100111010111000111100001100010011001100101110001111000011000110011011000111010010111000111100000110001011000010111111001011100011110000011000001100010011100110101110001111000001110000011100100100111;
			-9: data_out = 0110001000100111010111000111100001100010011001100101110001111000011000110011010001011100011110000011000000110110010111000111100000110000011000100110011101011100011110000110000100111000010100110111010100100111;
			-8: data_out = 0110001000100111010111000111100001100010011001100101110001111000011000110011000101011100011110000110010000110000011011000101110001111000001110010011011001011100011110000011100001100100010111000111100000111001011001010101110001111000001100010011100100100111;
			-7: data_out = 0110001000100111010111000111100001100010011001100101110001111000011000100110011000110010010111000111100001100100001101000100110001001111011000100101110001111000011001000011001100100111;
			-6: data_out = 0110001000100111010111000111100001100010011001100101110001111000011000100110000101011100011110000110001100110010011000000101110001111000001110010110001000111100010101110110101100100111;
			-5: data_out = 0110001000100111010111000111100001100010011001100101110001111000011000100011011001001111010111000111100001100100001101100101110001111000011000100011100001011100011110000110001100110010010111000111100000111000001100010101110001111000001100000011001000100111;
			-4: data_out = 0110001000100111010111000111100001100010011001100101110001111000011000100011000101011100011110000110010001100010010111000111100000111000011001100110110101101010010100010010100000100111;
			-3: data_out = 011000100010011101011100011110000110001001100110010111000111100001100001011000010101110001111000011000110110001001011100011110000110001100110111010010000101110001111000011001010110011001011100011110000110001100111001010111000111001000100111;
			-2: data_out = 0110001000100010010111000111100001100010011001100101110001111000011000010011000101011100011110000110010001100101010110000101110001111000011000110011100101011100011110000110011000110111010111000111100001100100011000110010011100100010;
			-1: data_out = 0110001000100111010111000111100001100010011001100101110001111000001110010011000101011100011110000110010001100110010111000111100000110000011000100010101101011100011110000011100000111001010111000111100001100100011001000101110001111000001100010110010100100111;
			0: data_out = 0110001000100111010111000111100000110000001100000101110001111000001100000011000001011100011110000011000000110000010111000111100000110000001100000101110001111000001100000011000001011100011110000011000000110000010111000111100000110000001100000101110001111000001100000011000000100111;
			1: data_out = 0110001000100111001111110101110001111000001110010011000101011100011110000110010001100110010111000111100000110000011000100010101101011100011110000011100000111001010111000111100001100100011001000101110001111000001100010110010100100111;
			2: data_out = 0110001000100010001111110101110001111000011000010011000101011100011110000110010001100101010110000101110001111000011000110011100101011100011110000110011000110111010111000111100001100100011000110010011100100010;
			3: data_out = 011000100010011100111111010111000111100001100001011000010101110001111000011000110110001001011100011110000110001100110111010010000101110001111000011001010110011001011100011110000110001100111001010111000111001000100111;
			4: data_out = 0110001000100111001111110101110001111000011000100011000101011100011110000110010001100010010111000111100000111000011001100110110101101010010100010010100000100111;
			5: data_out = 0110001000100111001111110101110001111000011000100011011001001111010111000111100001100100001101100101110001111000011000100011100001011100011110000110001100110010010111000111100000111000001100010101110001111000001100000011001000100111;
			6: data_out = 0110001000100111001111110101110001111000011000100110000101011100011110000110001100110010011000000101110001111000001110010110001000111100010101110110101100100111;
			7: data_out = 0110001000100111001111110101110001111000011000100110011000110010010111000111100001100100001101000100110001001111011000100101110001111000011001000011001100100111;
			8: data_out = 0110001000100111001111110101110001111000011000110011000101011100011110000110010000110000011011000101110001111000001110010011011001011100011110000011100001100100010111000111100000111001011001010101110001111000001100010011100100100111;
			9: data_out = 0110001000100111001111110101110001111000011000110011010001011100011110000011000000110110010111000111100000110000011000100110011101011100011110000110000100111000010100110111010100100111;
			10: data_out = 0110001000100111001111110101110001111000011000110011011000111010010111000111100000110001011000010111111001011100011110000011000001100010011100110101110001111000001110000011100100100111;
			11: data_out = 0110001000100111001111110101110001111000011000110011100001101100011011010101110001111000011001000110010001110110011000100100111100100111;
			12: data_out = 0110001000100111001111110101110001111000011000110110000101011100011110000011100101100011010111000111100001100100001110010101110001111000011000010110001101000010010110000101110001111000011001100011010100100111;
			13: data_out = 0110001000100111001111110101110001111000011000110110001101011100011110000110001101100010001100100011011001011100011110000110001101100100010111000111100001100011001101100111010100100111;
			14: data_out = 0110001000100111001111110101110001111000011000110110010101011100011110000110011000110111010010110101110001111000011001100011001001011100011110000110010100110100010111000111100001100010001110010101110001111000001100010110010000100111;
			15: data_out = 0110001000100111001111110101110001111000011001000011000001011100011110000011100100110000011111010101110001111000011000110011000101011100011110000011100100110011010111000111100000110000001101100101110001111000001110010011000000100111;
			16: data_out = 011000100010011100111111010111000111100001100100001100010101110001111000011000010011010001011100011011100101110001111000011001000110010000110010010111000111100000111000011001010010100100100111;
			17: data_out = 0110001000100111001111110101110001111000011001000011001001011100011110000110001000110110001101110101110001111000011000110110011001011100011110000011100000110011010111000111100001100100001101010101110001111000011000110011100000100111;
			18: data_out = 0110001000100111001111110101110001111000011001000011001101011100011110000110001100110110010111000111100001100101011001100011011100101111010111000111100001100101001110010100111100100111;
			19: data_out = 0110001000100111001111110101110001111000011001000011010001011100011110000110010000110110010111000111100000110001011000100101110001111000011001000011000001011100011110000011000000110000010111000111100001100011011001000101110001111000011001000110001000100111;
			20: data_out = 0110001000100111001111110101110001111000011001000011010101011100011110000110010100110011010111000111100001100001001110000111010001011100011110000011100001100001010111000111100000110000011000100101110001111000011001100011010100100111;
			21: data_out = 0110001000100111001111110101110001111000011001000011011001011100011110000110010101100110010111000111100000111000001100000101110001111000001100010110011001011100011110000110001101100101010111000111100001100100001100110011110000100111;
			22: data_out = 0110001000100111001111110101110001111000011001000011011101011100011110000110011000111001010111000111100000111000011001000101110001111000011001010110010101011100011110000110010100110101010111000111100000111001001101100101110001111000001110000011000100100111;
			23: data_out = 0110001000100111001111110101110001111000011001000011100101011100011110000011000000110001010111000111100001100010011001000010001001011100011110000011100100111000010111000111100001100110011001100101110001111000011000010110000100100111;
			24: data_out = 0110001000100111001111110101110001111000011001000110000101011100011110000011000000110111010111000111100001100110001110010010000101011100011110000011000000110110010111000111100000110001011000010101110001111000011001000011000000100111;
			25: data_out = 0110001000100111001111110101110001111000011001000110001001011100011110000011000001100011001011010111011100110111010111000111100000111001001110000101001100100111;
			26: data_out = 0110001000100111001111110101110001111000011001000110001101011100011110000011000001100101010001010101110001111000011001000110000101011100011110000110001001100101010111000111100000110000001101010101110001111000011000110011100000100111;
			27: data_out = 0110001000100111001111110101110001111000011001000110010001011100011110000011000001100101001011100010101101000100010111000111100001100100011001010101110001111000001100000011000000100111;
			28: data_out = 0110001000100111001111110101110001111000011001000110010101011100011110000011000001100010010111000111100001100100001100100111010000100100010100000111100100100111;
			29: data_out = 0110001000100111001111110101110001111000011001000110011001011100011110000011000000110111010111000111100000110001011001010101110001111000011001010110010001011100011110000110010101100110010111000111100001100001001100000101110001111000011001010110010000100111;
			30: data_out = 0110001000100111001111110101110001111000011001000110011001011100011110000110011001100110010111000111100001100110011001100101110001111000011001100110011001011100011110000110011001100110010111000111100001100110011001100101110001111000011001100110011000100111;
			31: data_out = 0110001000100111001111110101110001111000011001010011000001111011001100010010000001011100011110000110011001100100010111000111100001100100011001100101110001111000001100010011001100100111;
			32: data_out = 0110001000100111001111110101110001111000011001010011000001011100011110000110011000110101010111000111100000110001001110010011111001011100011110000110000101100011010111000111100001100100011001000010101000100111;
			33: data_out = 0110001000100111001111110101110001111000011001010011000101101101010111000111100001100001011001010101110001111000011001000011011101110000011101110101110001111000001100010110010000100111;
			34: data_out = 0110001000100111001111110101110001111000011001010011000101011100011110000110010100110100010111000111100001100101001110000101110001111000001110000011010001011100011110000011000100110001010111000111100001100110011001000101110001111000001100010011001100100111;
			35: data_out = 0110001000100111001111110101110001111000011001010011001001011010010111000111100001100010011000110101110001111000011001100011100001111100010010010111100000100111;
			36: data_out = 0110001000100111001111110101110001111000011001010011001001011100011110000110001101100110001000110101110001111000001100000011010001110101010110100101111000100111;
			37: data_out = 0110001000100111001111110101110001111000011001010011001101000010010111000111100000110001001100010101110001111000001110010011010001010101010111000111100001100010011001010101110001111000011000100011011000100111;
			38: data_out = 0110001000100111001111110101110001111000011001010011001101011100011110000110001000110011010111000111100000110111011001100101110001111000011000100011000101011100011110000110001001100100010111000111100001100011001110010011100000100111;
			39: data_out = 0110001000100111001111110101110001111000011001010011010000100011011001000101110001111000001110000011010001001000011110100101110001111000011000100110010000100111;
			40: data_out = 0110001000100111001111110101110001111000011001010011010001011100011110000011100100110001010111000111100001100010001101110101001000111100010111000111100000110001001101100101110001111000001100010110001100100111;
			41: data_out = 0110001000100111001111110101110001111000011001010011010001011100011110000110011001100101011011110101110001111000001110000011000100111000010011110101110001111000011001000011001100100111;
			42: data_out = 0110001000100111001111110101110001111000011001010011010101101001010111000111100000111000001101000101110001111000001110010011011001011100011110000110010100110010010111000111100000110000011000100101110001111000011001000011100000100111;
			43: data_out = 0110001000100111001111110101110001111000011001010011010101011100011110000110010000110010010111000111100001100101011001010011100101011100011110000011100001100011010111000111100000111001011000110010101100100111;
			44: data_out = 0110001000100111001111110101110001111000011001010011011000111010010111000111100001100001001101000011000001011100011110000110010100110000011100110101110001111000001100010011000000100111;
			45: data_out = 0110001000100111001111110101110001111000011001010011011001011100011110000110000100110000010111000111100000111001011001010110011001011100011110000011011101100110001110110101110001111000011000110110001100100111;
			46: data_out = 0110001000100111001111110101110001111000011001010011011101011100011110000011000000110100010111000111100001100100001101000101110001111000011001010011011001011100011110000110000100110101010011010011100000100111;
			47: data_out = 0110001000100111001111110101110001111000011001010011011101100111001111110101110001111000011001010011000001011100011110000110001100111000011010010101110001111000001110000011001000100111;
			48: data_out = 0110001000100111001111110101110001111000011001010011011101011100011110000110001100110111010111000111100001100100001101110101110001111000011000010011100000110011010111000111100001100010011001010101110001111000011000110011000100100111;
			49: data_out = 0110001000100111001111110101110001111000011001010011100000100110010111000111100000111001001101000101110001111000011000100011010001011100011110000110000100110001010111000111100000110001011000110011011100100111;
			50: data_out = 0110001000100111001111110101110001111000011001010011100001011100011110000011100000110011011011110101110001111000011000010011001001011100011110000110001101100110010100000011100100100111;
			51: data_out = 0110001000100010001111110101110001111000011001010011100001011100011110000110010001100101011000010011010101011100011110000011000100110101010111000111100001100001001100110010011100100010;
			52: data_out = 0110001000100111001111110101110001111000011001010011100100110111011000100101001101011100011110000110011000110100011000110101110001111000011001000011001000100111;
			53: data_out = 0110001000100111001111110101110001111000011001010011100101011100011110000011100001100101011011000101110001111000001100000110010101011100011110000110000100110010011110100101110001111000001100010011010000100111;
			54: data_out = 0110001000100111001111110101110001111000011001010011100101011100011110000110010100110011011101110101110001111000001110010110001001011100011110000011100100110111010111000111100001100110001101000101110001111000011000010011100000100111;
			55: data_out = 0110001000100111001111110101110001111000011001010110000100110110011111100101100101011100011110000011000100110101010111000111100000111000001101110100011100100111;
			56: data_out = 0110001000100111001111110101110001111000011001010110000101011100011110000011100000110111011110010101110001111000011000110110010001011100011110000110000100111000010111000111100001100101011001010101110001111000011000010011010100100111;
			57: data_out = 0110001000100111001111110101110001111000011001010110000101011100011110000110010000110110011000110101110001111000011000010011100001011100011110000110000101100101001011110101110001111000011001000110001000100111;
			58: data_out = 0110001000100111001111110101110001111000011001010110001000100011001101010101110001111000011000110011001001011100011110000110001101100100010111000111100001100001001110010100010100100111;
			59: data_out = 0110001000100111001111110101110001111000011001010110001001101101010111000111100001100101011000010101110001111000001100010110010101110110010111000111100001100101011000010101110001111000011001000110010000100111;
			60: data_out = 0110001000100111001111110101110001111000011001010110001001011100011110000110001000110110011110100101110001111000011001010011100001011000010011000101110001111000011000010110000100100111;
			61: data_out = 0110001000100111001111110101110001111000011001010110001001011100011110000110011001100011010111000111100001100101001100100111011101011100011110000110010000110011001110010101110001111000011000110011011000100111;
			62: data_out = 0110001000100010001111110101110001111000011001010110001101000001010111000111100000110001011000100100111101101101001001110101110001111000001100000011011100100010;
			63: data_out = 0110001000100111001111110101110001111000011001010110001101011100011110000011100000110011001000000101110001111000001100010110010000111101001011000110110000100111;
			64: data_out = 0110001000100111001111110101110001111000011001010110001101011100011110000110001100110010010111000111100001100101011000100101110001111000011000100110001001010110001110000101110001111000011000110110000100100111;
			65: data_out = 0110001000100111001111110101110001111000011001010110010001011100011110000011000000110000011110010011000000101101010111000111100001100100001101110110011100100111;
			66: data_out = 0110001000100111001111110101110001111000011001010110010000111011010111000111100001100011001100110101110001111000011000010110010101011100011110000110011001100110010111000111100000110111011001100101110001111000001110010011010100100111;
			67: data_out = 0110001000100111001111110101110001111000011001010110010001110100010111000111100001100011001101100101110001111000001110010011100000101100011001100110111000100111;
			68: data_out = 0110001000100111001111110101110001111000011001010110010001011100011110000110000101100010011111010111100101011100011110000011100100110111010111000111100001100011011000100101100000100111;
			69: data_out = 0110001000100111001111110101110001111000011001010110010001011100011110000110010001100110010111000111100001100101001101000101110001111000001100000110010101011100011110000110011001100110010111000111100001100010001110000101110001111000001100000011010100100111;
			70: data_out = 0110001000100111001111110101110001111000011001010110010101011100011110000011000100110001010111000111100001100110001101100100001001010010001011010101110001111000001100010110001000100111;
			71: data_out = 0110001000100111001111110101110001111000011001010110010101000001010111000111100001100010001100000010101101011100011110000110011001100101010111000111100001100010001101000101110001111000011000110110000100100111;
			72: data_out = 0110001000100111001111110101110001111000011001010110010101101111010111000111100000110000011001010101110001111000001100010011001101000100010101000101110001111000011001100110011000100111;
			73: data_out = 0110001000100111001111110101110001111000011001010110010101011100011110000011100101100001010111000111100000110000011000110110111001111011010111000111100001100100011000100101110001111000001100010110011000100111;
			74: data_out = 0110001000100111001111110101110001111000011001010110010101011100011110000110001100110010010111000111100001100001001101110101110001111000011001010011001101011110011110110101110001111000001110000011000000100111;
			75: data_out = 0110001000100111001111110101110001111000011001010110010101011100011110000110010100111000010111000111100001100100011001000100011101001000010111000111100001100010011001100101110001111000001100010011010100100111;
			76: data_out = 0110001000100111001111110101110001111000011001010110011001011100011110000011000001100011010111000111100001100001001110010101110001111000001110010110011001111001010111000111100001100010011000010010010100100111;
			77: data_out = 011000100010011100111111010111000111100001100101011001100010111001011100011011100010000101001110010111000111100000111000001101110101110001111000001100000110011000100111;
			78: data_out = 0110001000100111001111110101110001111000011001010110011001001100010111000111100001100110011000110011001001111010010111000111100000110000001100000101110001111000001101110110011000100111;
			79: data_out = 0110001000100111001111110101110001111000011001010110011001101001011111010110100100111000010111000111100001100010001101100101110001111000011000110011001000100111;
			80: data_out = 0110001000100111001111110101110001111000011001010110011001011100011110000011100000110011010111000111100000111000011000100101110001111000001110000110001101011100011110000011100000110001010111000111100000110001011000110101110001111000001100010011011100100111;
			81: data_out = 011000100010011100111111010111000111100001100101011001100101110001111000001110010110001000100100010111000111100000111001001101000010111101011100011110000110010100110100010111000101110000100111;
			82: data_out = 0110001000100111001111110101110001111000011001010110011001011100011110000110001000110000010001100101110001111000011000010011100100110000010111000111100000111001001101000111100100100111;
			83: data_out = 0110001000100111001111110101110001111000011001010110011001011100011110000110001100110010010111000111100001100110001100000010010101011100011110000110000100110010001111100101110001111000001110000110001000100111;
			84: data_out = 0110001000100111001111110101110001111000011001010110011001011100011110000110010000110011010111000111100000110001011001100101110001111000001110010011010001011100011110000110011000111000011001110101110001111000011000110011011000100111;
