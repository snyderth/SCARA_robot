module degrees_to_steps(input 	signed [31:0] dtheta1,
								input 	signed [31:0] dtheta2,
								output 	logic dir1,
								output 	logic dir2,
								output 	logic [7:0] steps1,
								output	logic [7:0] steps2);
								
			
								
								
								
endmodule
								