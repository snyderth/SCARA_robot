module ScaraController();



endmodule
