/***************************************************
*	File: 		CosDeg
*	Author: 		Thomas Snyder
*	Date:			2/5/2020
*	Description:Cosine Function inputing a signed integer
*					in degrees and outputing a double
					precision floating point number.
*	Parameters:
*				None
*	Dependencies:
*				None
*
***************************************************/
module	CosDeg(input	signed	[8:0]	data_in,
			output logic [63:0] data_out);


	always_comb
		case(data_in)
			 -180: data_out = 64'b1011111111110000000000000000000000000000000000000000000000000000;

			 -179: data_out = 64'b1011111111101111111111101100000010010111111011010001111101110111;

			 -178: data_out = 64'b1011111111101111111110110000001001111000101011011111111001101001;

			 -177: data_out = 64'b1011111111101111111101001100010111101100111110011000001000000011;

			 -176: data_out = 64'b1011111111101111111011000000101101110001010011110101100100110000;

			 -175: data_out = 64'b1011111111101111111000001101001110110011111011100100011100111110;

			 -174: data_out = 64'b1011111111101111110100110001111110010100110001101000110101101110;

			 -173: data_out = 64'b1011111111101111110000101111000000100101011010000111010001111101;

			 -172: data_out = 64'b1011111111101111101100000100011010101000111011101111011110000110;

			 -171: data_out = 64'b1011111111101111100110110010010010010011111001101001000111100010;

			 -170: data_out = 64'b1011111111101111100000111000101110001100001100000011001000000001;

			 -169: data_out = 64'b1011111111101111011010010111110101101000111000000101001101111011;

			 -168: data_out = 64'b1011111111101111010011001111110000110010000110100100001011111001;

			 -167: data_out = 64'b1011111111101111001011100000101000100000111001111000111010110100;

			 -166: data_out = 64'b1011111111101111000011001010100110011111000010111010011011011100;

			 -165: data_out = 64'b1011111111101110111010001101110101000110110100111011000100110101;

			 -164: data_out = 64'b1011111111101110110000101010011111100010111000101001001111010100;

			 -163: data_out = 64'b1011111111101110100110100000110001101101111110010011101011011100;

			 -162: data_out = 64'b1011111111101110011011110000111000010010101110110001110111000000;

			 -161: data_out = 64'b1011111111101110010000011011000000101011011011110000100010001110;

			 -160: data_out = 64'b1011111111101110000100011111011001000001101111000010111000111110;

			 -159: data_out = 64'b1011111111101101110111111110010000001110011000111000100100111101;

			 -158: data_out = 64'b1011111111101101101010110111110101111000111101011000111110110001;

			 -157: data_out = 64'b1011111111101101011101001100011010010111100001000100000101000101;

			 -156: data_out = 64'b1011111111101101001110111100001110101110010100011001010010010001;

			 -155: data_out = 64'b1011111111101101000000000111100100101111011110100100101001111000;

			 -154: data_out = 64'b1011111111101100110000101110101110111010100111010010111000100001;

			 -153: data_out = 64'b1011111111101100100000110010000000011100011111101100100001111110;

			 -152: data_out = 64'b1011111111101100010000010001101101001110101010011000111001111110;

			 -151: data_out = 64'b1011111111101011111111001110001001110111000010101001000110000011;

			 -150: data_out = 64'b1011111111101011101101100111101011100111100010101011100110111111;

			 -149: data_out = 64'b1011111111101011011011011110101000011101101001001001001010000111;

			 -148: data_out = 64'b1011111111101011001000110011010111000001111101101011000011101010;

			 -147: data_out = 64'b1011111111101010110101100110001110100111110100101011110100000101;

			 -146: data_out = 64'b1011111111101010100001110111100111001100110010010010011011110110;

			 -145: data_out = 64'b1011111111101010001101100111111001011000001100011001000010000101;

			 -144: data_out = 64'b1011111111101001111000110111011110011010101011111111010010101010;

			 -143: data_out = 64'b1011111111101001100011100110110000001101101101101001011011000010;

			 -142: data_out = 64'b1011111111101001001101110110001001010011000001001100001100011101;

			 -141: data_out = 64'b1011111111101000110111100110000100110100001000100110101100010000;

			 -140: data_out = 64'b1011111111101000100000110110111110100001110110001010011011000001;

			 -139: data_out = 64'b1011111111101000001001101001010010110011101001110010011101011010;

			 -138: data_out = 64'b1011111111100111110001111101011110100111001101101010010001111001;

			 -137: data_out = 64'b1011111111100111011001110011111111011111110010000100111110111111;

			 -136: data_out = 64'b1011111111100111000001001101010011100101101000100101100111011110;

			 -135: data_out = 64'b1011111111100110101000001001111001100101011110011001010010101010;

			 -134: data_out = 64'b1011111111100110001110101010010000101111110110000011110111011100;

			 -133: data_out = 64'b1011111111100101110100101110111000111000100000011111111010000110;

			 -132: data_out = 64'b1011111111100101011010011000010010010101110101010010101101000011;

			 -131: data_out = 64'b1011111111100100111111100110111110000000001010010101000110100101;

			 -130: data_out = 64'b1011111111100100100100011011011101010001001010110001111110001010;

			 -129: data_out = 64'b1011111111100100001000110110010010000011001101011011000011001110;

			 -128: data_out = 64'b1011111111100011101100110111111110110000101010010101000011000100;

			 -127: data_out = 64'b1011111111100011010000100001000110010011001111111011110001100000;

			 -126: data_out = 64'b1011111111100010110011110010001100000011010111011111001010001110;

			 -125: data_out = 64'b1011111111100010010110101011110011110111011000111010000001100001;

			 -124: data_out = 64'b1011111111100001111001001110100010000010111110000011011010100011;

			 -123: data_out = 64'b1011111111100001011011011010111011010110010101011011011100000001;

			 -122: data_out = 64'b1011111111100000111101010001100100111101100100010100011011000101;

			 -121: data_out = 64'b1011111111100000011110110011000100011111111000011001010101111101;

			 -120: data_out = 64'b1011111111011111111111111111111111111101110001100100110000000001;

			 -119: data_out = 64'b1011111111011111000001110001111011101011101101010001000011111111;

			 -118: data_out = 64'b1011111111011110000010111101001001110001111010010010100011100010;

			 -117: data_out = 64'b1011111111011101000011100010111000101001000010010110001001001010;

			 -116: data_out = 64'b1011111111011100000011100100010111011000100000100111100010111111;

			 -115: data_out = 64'b1011111111011011000011000010110101110100111111000011110000000011;

			 -114: data_out = 64'b1011111111011010000001111111100100011110110010110011000001111011;

			 -113: data_out = 64'b1011111111011001000000011011110100100000010111101100011111000001;

			 -112: data_out = 64'b1011111111010111111110011000110111101100101011000101000010011010;

			 -111: data_out = 64'b1011111111010110111011111000000000011101100101101011111000011010;

			 -110: data_out = 64'b1011111111010101111000111010100001110010010100110110010101101111;

			 -109: data_out = 64'b1011111111010100110101100001101111001101110010111101001011100110;

			 -108: data_out = 64'b1011111111010011110001101110111100110100111111001101010111101011;

			 -107: data_out = 64'b1011111111010010101101100011011111001101010100101110010011111101;

			 -106: data_out = 64'b1011111111010001101001000000101011011011000000111111101000010001;

			 -105: data_out = 64'b1011111111010000100100000111110110111111011001110000100000110101;

			 -104: data_out = 64'b1011111111001110111101110100101111101110100100100101011111101010;

			 -103: data_out = 64'b1011111111001100110010110011001000110010100000010110111011001001;

			 -102: data_out = 64'b1011111111001010100111001101100110100111111111000111011010100000;

			 -101: data_out = 64'b1011111111001000011011000110110111011001001101110101111100000011;

			 -100: data_out = 64'b1011111111000110001110100001101001111001110100111011011010110101;

			 -99: data_out = 64'b1011111111000100000001100000101101100011011110000100001001010110;

			 -98: data_out = 64'b1011111111000001110100000110110010010010011001011001101110100100;

			 -97: data_out = 64'b1011111110111111001100101101010001000100000100000011110001010011;

			 -96: data_out = 64'b1011111110111010110000100110000010010011000011101100101111101000;

			 -95: data_out = 64'b1011111110110110010011111101011010110000101001110100100000110111;

			 -94: data_out = 64'b1011111110110001110110111000111101100101011000100001110111101101;

			 -93: data_out = 64'b1011111110101010110010111100011100111001000001101100100111011101;

			 -92: data_out = 64'b1011111110100001110111100101100010111010001101111001011000111011;

			 -91: data_out = 64'b1011111110010001110111110000101100001100010111010101010001001001;

			 -90: data_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;

			 -89: data_out = 64'b0011111110010001110111110000101101001010000001110000000001011000;

			 -88: data_out = 64'b0011111110100001110111100101100011011001000010001101000011111101;

			 -87: data_out = 64'b0011111110101010110010111100011101010111110100100000001000100101;

			 -86: data_out = 64'b0011111110110001110110111000111101110100110000111000010101110110;

			 -85: data_out = 64'b0011111110110110010011111101011011000000000000110100100000001100;

			 -84: data_out = 64'b0011111110111010110000100110000010100010011001000011000110001001;

			 -83: data_out = 64'b0011111110111111001100101101010001010011010111011101010110010111;

			 -82: data_out = 64'b0011111111000001110100000110110010011010000001111110100101011000;

			 -81: data_out = 64'b0011111111000100000001100000101101101011000101010111100010111110;

			 -80: data_out = 64'b0011111111000110001110100001101010000001011010110011110111001010;

			 -79: data_out = 64'b0011111111001000011011000110110111100000110010001001111100101111;

			 -78: data_out = 64'b0011111111001010100111001101100110101111100001101101100011011000;

			 -77: data_out = 64'b0011111111001100110010110011001000111010000001000101110010000110;

			 -76: data_out = 64'b0011111111001110111101110100101111110110000011010011101100111001;

			 -75: data_out = 64'b0011111111010000100100000111110111000011001000000010100111111000;

			 -74: data_out = 64'b0011111111010001101001000000101011011110101110001000000110100000;

			 -73: data_out = 64'b0011111111010010101101100011011111010001000000101000100001101000;

			 -72: data_out = 64'b0011111111010011110001101110111100111000101001110100101110010010;

			 -71: data_out = 64'b0011111111010100110101100001101111010001011100001101000110100001;

			 -70: data_out = 64'b0011111111010101111000111010100001110101111100101010010001110110;

			 -69: data_out = 64'b0011111111010110111011111000000000100001001011111111010100100010;

			 -68: data_out = 64'b0011111111010111111110011000110111110000001111110011011111001101;

			 -67: data_out = 64'b0011111111011001000000011011110100100011111010110001011111000110;

			 -66: data_out = 64'b0011111111011010000001111111100100100010010100001010001001111010;

			 -65: data_out = 64'b0011111111011011000011000010110101111000011110101000100110111000;

			 -64: data_out = 64'b0011111111011100000011100100010111011011111110010101110001101011;

			 -63: data_out = 64'b0011111111011101000011100010111000101100011110001001011011000110;

			 -62: data_out = 64'b0011111111011110000010111101001001110101010100000110100110011011;

			 -61: data_out = 64'b0011111111011111000001110001111011101111000101000001101000000101;

			 -60: data_out = 64'b0011111111100000000000000000000000000000100011100110110100000000;

			 -59: data_out = 64'b0011111111100000011110110011000100100001100010000111110110101100;

			 -58: data_out = 64'b0011111111100000111101010001100100111111001100111010111100101000;

			 -57: data_out = 64'b0011111111100001011011011010111011010111111100110111111011110111;

			 -56: data_out = 64'b0011111111100001111001001110100010000100100100010011110111101001;

			 -55: data_out = 64'b0011111111100010010110101011110011111000111101111100011100010010;

			 -54: data_out = 64'b0011111111100010110011110010001100000100111011010001100100100100;

			 -53: data_out = 64'b0011111111100011010000100001000110010100110010011100001110111000;

			 -52: data_out = 64'b0011111111100011101100110111111110110010001011100001101000101000;

			 -51: data_out = 64'b0011111111100100001000110110010010000100101101010001110111101101;

			 -50: data_out = 64'b0011111111100100100100011011011101010010101001010001001001111101;

			 -49: data_out = 64'b0011111111100100111111100110111110000001100111011010110011110010;

			 -48: data_out = 64'b0011111111100101011010011000010010010111010000111101000111100000;

			 -47: data_out = 64'b0011111111100101110100101110111000111001111010101101001111100000;

			 -46: data_out = 64'b0011111111100110001110101010010000110001001110110010010111001110;

			 -45: data_out = 64'b0011111111100110101000001001111001100110110101100111001110000100;

			 -44: data_out = 64'b0011111111100111000001001101010011100110111110010001010001101100;

			 -43: data_out = 64'b0011111111100111011001110011111111100001000110001100101101001010;

			 -42: data_out = 64'b0011111111100111110001111101011110101000100000001100011011000010;

			 -41: data_out = 64'b0011111111101000001001101001010010110100111010101101011010100001;

			 -40: data_out = 64'b0011111111101000100000110110111110100011000101011100100111001010;

			 -39: data_out = 64'b0011111111101000110111100110000100110101010110001110100100100011;

			 -38: data_out = 64'b0011111111101001001101110110001001010100001101001000010000000001;

			 -37: data_out = 64'b0011111111101001100011100110110000001110110111111000001011000101;

			 -36: data_out = 64'b0011111111101001111000110111011110011011110100011111010010100111;

			 -35: data_out = 64'b0011111111101010001101100111111001011001010011001000110111011111;

			 -34: data_out = 64'b0011111111101010100001110111100111001101110111010000101110011100;

			 -33: data_out = 64'b0011111111101010110101100110001110101000110111110111001101101111;

			 -32: data_out = 64'b0011111111101011001000110011010111000010111111000010010000101000;

			 -31: data_out = 64'b0011111111101011011011011110101000011110101000101010111000110110;

			 -30: data_out = 64'b0011111111101011101101100111101011101000100000010110101000001101;

			 -29: data_out = 64'b0011111111101011111111001110001001110111111110011100001100110100;

			 -28: data_out = 64'b0011111111101100010000010001101101001111100100010010111011101011;

			 -27: data_out = 64'b0011111111101100100000110010000000011101010111101100010110010111;

			 -26: data_out = 64'b0011111111101100110000101110101110111011011101010111011001101110;

			 -25: data_out = 64'b0011111111101101000000000111100100110000010010101100110100011010;

			 -24: data_out = 64'b0011111111101101001110111100001110101111000110100100000101000111;

			 -23: data_out = 64'b0011111111101101011101001100011010011000010001010000100001101001;

			 -22: data_out = 64'b0011111111101101101010110111110101111001101011100110001000111011;

			 -21: data_out = 64'b0011111111101101110111111110010000001111000101000101100011000100;

			 -20: data_out = 64'b0011111111101110000100011111011001000010011001001110110011110111;

			 -19: data_out = 64'b0011111111101110010000011011000000101100000011111010100101010001;

			 -18: data_out = 64'b0011111111101110011011110000111000010011010100111001010000000110;

			 -17: data_out = 64'b0011111111101110100110100000110001101110100010010111101011000010;

			 -16: data_out = 64'b0011111111101110110000101010011111100011011010101001001000011010;

			 -15: data_out = 64'b0011111111101110111010001101110101000111010100110110001101000000;

			 -14: data_out = 64'b0011111111101111000011001010100110011111100000110000001010110110;

			 -13: data_out = 64'b0011111111101111001011100000101000100001010101101000101100010000;

			 -12: data_out = 64'b0011111111101111010011001111110000110010100000001101011100101110;

			 -11: data_out = 64'b0011111111101111011010010111110101101001001111100111011110001010;

			 -10: data_out = 64'b0011111111101111100000111000101110001100100001011101111010010001;

			 -9: data_out = 64'b0011111111101111100110110010010010010100001100111100000001000111;

			 -8: data_out = 64'b0011111111101111101100000100011010101001001100111010000110111010;

			 -7: data_out = 64'b0011111111101111110000101111000000100101101001001001010100100110;

			 -6: data_out = 64'b0011111111101111110100110001111110010100111110100001111111011011;

			 -5: data_out = 64'b0011111111101111111000001101001110110100000110010100011101101010;

			 -4: data_out = 64'b0011111111101111111011000000101101110001011100011100001111000001;

			 -3: data_out = 64'b0011111111101111111101001100010111101101000100110101010001001001;

			 -2: data_out = 64'b0011111111101111111110110000001001111000101111110011011001100001;

			 -1: data_out = 64'b0011111111101111111111101100000010010111111101011011101111001001;

			 0: data_out = 64'b0011111111110000000000000000000000000000000000000000000000000000;

			 1: data_out = 64'b0011111111101111111111101100000010010111111101011011101111001001;

			 2: data_out = 64'b0011111111101111111110110000001001111000101111110011011001100001;

			 3: data_out = 64'b0011111111101111111101001100010111101101000100110101010001001001;

			 4: data_out = 64'b0011111111101111111011000000101101110001011100011100001111000001;

			 5: data_out = 64'b0011111111101111111000001101001110110100000110010100011101101010;

			 6: data_out = 64'b0011111111101111110100110001111110010100111110100001111111011011;

			 7: data_out = 64'b0011111111101111110000101111000000100101101001001001010100100110;

			 8: data_out = 64'b0011111111101111101100000100011010101001001100111010000110111010;

			 9: data_out = 64'b0011111111101111100110110010010010010100001100111100000001000111;

			 10: data_out = 64'b0011111111101111100000111000101110001100100001011101111010010001;

			 11: data_out = 64'b0011111111101111011010010111110101101001001111100111011110001010;

			 12: data_out = 64'b0011111111101111010011001111110000110010100000001101011100101110;

			 13: data_out = 64'b0011111111101111001011100000101000100001010101101000101100010000;

			 14: data_out = 64'b0011111111101111000011001010100110011111100000110000001010110110;

			 15: data_out = 64'b0011111111101110111010001101110101000111010100110110001101000000;

			 16: data_out = 64'b0011111111101110110000101010011111100011011010101001001000011010;

			 17: data_out = 64'b0011111111101110100110100000110001101110100010010111101011000010;

			 18: data_out = 64'b0011111111101110011011110000111000010011010100111001010000000110;

			 19: data_out = 64'b0011111111101110010000011011000000101100000011111010100101010001;

			 20: data_out = 64'b0011111111101110000100011111011001000010011001001110110011110111;

			 21: data_out = 64'b0011111111101101110111111110010000001111000101000101100011000100;

			 22: data_out = 64'b0011111111101101101010110111110101111001101011100110001000111011;

			 23: data_out = 64'b0011111111101101011101001100011010011000010001010000100001101001;

			 24: data_out = 64'b0011111111101101001110111100001110101111000110100100000101000111;

			 25: data_out = 64'b0011111111101101000000000111100100110000010010101100110100011010;

			 26: data_out = 64'b0011111111101100110000101110101110111011011101010111011001101110;

			 27: data_out = 64'b0011111111101100100000110010000000011101010111101100010110010111;

			 28: data_out = 64'b0011111111101100010000010001101101001111100100010010111011101011;

			 29: data_out = 64'b0011111111101011111111001110001001110111111110011100001100110100;

			 30: data_out = 64'b0011111111101011101101100111101011101000100000010110101000001101;

			 31: data_out = 64'b0011111111101011011011011110101000011110101000101010111000110110;

			 32: data_out = 64'b0011111111101011001000110011010111000010111111000010010000101000;

			 33: data_out = 64'b0011111111101010110101100110001110101000110111110111001101101111;

			 34: data_out = 64'b0011111111101010100001110111100111001101110111010000101110011100;

			 35: data_out = 64'b0011111111101010001101100111111001011001010011001000110111011111;

			 36: data_out = 64'b0011111111101001111000110111011110011011110100011111010010100111;

			 37: data_out = 64'b0011111111101001100011100110110000001110110111111000001011000101;

			 38: data_out = 64'b0011111111101001001101110110001001010100001101001000010000000001;

			 39: data_out = 64'b0011111111101000110111100110000100110101010110001110100100100011;

			 40: data_out = 64'b0011111111101000100000110110111110100011000101011100100111001010;

			 41: data_out = 64'b0011111111101000001001101001010010110100111010101101011010100001;

			 42: data_out = 64'b0011111111100111110001111101011110101000100000001100011011000010;

			 43: data_out = 64'b0011111111100111011001110011111111100001000110001100101101001010;

			 44: data_out = 64'b0011111111100111000001001101010011100110111110010001010001101100;

			 45: data_out = 64'b0011111111100110101000001001111001100110110101100111001110000100;

			 46: data_out = 64'b0011111111100110001110101010010000110001001110110010010111001110;

			 47: data_out = 64'b0011111111100101110100101110111000111001111010101101001111100000;

			 48: data_out = 64'b0011111111100101011010011000010010010111010000111101000111100000;

			 49: data_out = 64'b0011111111100100111111100110111110000001100111011010110011110010;

			 50: data_out = 64'b0011111111100100100100011011011101010010101001010001001001111101;

			 51: data_out = 64'b0011111111100100001000110110010010000100101101010001110111101101;

			 52: data_out = 64'b0011111111100011101100110111111110110010001011100001101000101000;

			 53: data_out = 64'b0011111111100011010000100001000110010100110010011100001110111000;

			 54: data_out = 64'b0011111111100010110011110010001100000100111011010001100100100100;

			 55: data_out = 64'b0011111111100010010110101011110011111000111101111100011100010010;

			 56: data_out = 64'b0011111111100001111001001110100010000100100100010011110111101001;

			 57: data_out = 64'b0011111111100001011011011010111011010111111100110111111011110111;

			 58: data_out = 64'b0011111111100000111101010001100100111111001100111010111100101000;

			 59: data_out = 64'b0011111111100000011110110011000100100001100010000111110110101100;

			 60: data_out = 64'b0011111111100000000000000000000000000000100011100110110100000000;

			 61: data_out = 64'b0011111111011111000001110001111011101111000101000001101000000101;

			 62: data_out = 64'b0011111111011110000010111101001001110101010100000110100110011011;

			 63: data_out = 64'b0011111111011101000011100010111000101100011110001001011011000110;

			 64: data_out = 64'b0011111111011100000011100100010111011011111110010101110001101011;

			 65: data_out = 64'b0011111111011011000011000010110101111000011110101000100110111000;

			 66: data_out = 64'b0011111111011010000001111111100100100010010100001010001001111010;

			 67: data_out = 64'b0011111111011001000000011011110100100011111010110001011111000110;

			 68: data_out = 64'b0011111111010111111110011000110111110000001111110011011111001101;

			 69: data_out = 64'b0011111111010110111011111000000000100001001011111111010100100010;

			 70: data_out = 64'b0011111111010101111000111010100001110101111100101010010001110110;

			 71: data_out = 64'b0011111111010100110101100001101111010001011100001101000110100001;

			 72: data_out = 64'b0011111111010011110001101110111100111000101001110100101110010010;

			 73: data_out = 64'b0011111111010010101101100011011111010001000000101000100001101000;

			 74: data_out = 64'b0011111111010001101001000000101011011110101110001000000110100000;

			 75: data_out = 64'b0011111111010000100100000111110111000011001000000010100111111000;

			 76: data_out = 64'b0011111111001110111101110100101111110110000011010011101100111001;

			 77: data_out = 64'b0011111111001100110010110011001000111010000001000101110010000110;

			 78: data_out = 64'b0011111111001010100111001101100110101111100001101101100011011000;

			 79: data_out = 64'b0011111111001000011011000110110111100000110010001001111100101111;

			 80: data_out = 64'b0011111111000110001110100001101010000001011010110011110111001010;

			 81: data_out = 64'b0011111111000100000001100000101101101011000101010111100010111110;

			 82: data_out = 64'b0011111111000001110100000110110010011010000001111110100101011000;

			 83: data_out = 64'b0011111110111111001100101101010001010011010111011101010110010111;

			 84: data_out = 64'b0011111110111010110000100110000010100010011001000011000110001001;

			 85: data_out = 64'b0011111110110110010011111101011011000000000000110100100000001100;

			 86: data_out = 64'b0011111110110001110110111000111101110100110000111000010101110110;

			 87: data_out = 64'b0011111110101010110010111100011101010111110100100000001000100101;

			 88: data_out = 64'b0011111110100001110111100101100011011001000010001101000011111101;

			 89: data_out = 64'b0011111110010001110111110000101101001010000001110000000001011000;

			 90: data_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;

			 91: data_out = 64'b1011111110010001110111110000101100001100010111010101010001001001;

			 92: data_out = 64'b1011111110100001110111100101100010111010001101111001011000111011;

			 93: data_out = 64'b1011111110101010110010111100011100111001000001101100100111011101;

			 94: data_out = 64'b1011111110110001110110111000111101100101011000100001110111101101;

			 95: data_out = 64'b1011111110110110010011111101011010110000101001110100100000110111;

			 96: data_out = 64'b1011111110111010110000100110000010010011000011101100101111101000;

			 97: data_out = 64'b1011111110111111001100101101010001000100000100000011110001010011;

			 98: data_out = 64'b1011111111000001110100000110110010010010011001011001101110100100;

			 99: data_out = 64'b1011111111000100000001100000101101100011011110000100001001010110;

			 100: data_out = 64'b1011111111000110001110100001101001111001110100111011011010110101;

			 101: data_out = 64'b1011111111001000011011000110110111011001001101110101111100000011;

			 102: data_out = 64'b1011111111001010100111001101100110100111111111000111011010100000;

			 103: data_out = 64'b1011111111001100110010110011001000110010100000010110111011001001;

			 104: data_out = 64'b1011111111001110111101110100101111101110100100100101011111101010;

			 105: data_out = 64'b1011111111010000100100000111110110111111011001110000100000110101;

			 106: data_out = 64'b1011111111010001101001000000101011011011000000111111101000010001;

			 107: data_out = 64'b1011111111010010101101100011011111001101010100101110010011111101;

			 108: data_out = 64'b1011111111010011110001101110111100110100111111001101010111101011;

			 109: data_out = 64'b1011111111010100110101100001101111001101110010111101001011100110;

			 110: data_out = 64'b1011111111010101111000111010100001110010010100110110010101101111;

			 111: data_out = 64'b1011111111010110111011111000000000011101100101101011111000011010;

			 112: data_out = 64'b1011111111010111111110011000110111101100101011000101000010011010;

			 113: data_out = 64'b1011111111011001000000011011110100100000010111101100011111000001;

			 114: data_out = 64'b1011111111011010000001111111100100011110110010110011000001111011;

			 115: data_out = 64'b1011111111011011000011000010110101110100111111000011110000000011;

			 116: data_out = 64'b1011111111011100000011100100010111011000100000100111100010111111;

			 117: data_out = 64'b1011111111011101000011100010111000101001000010010110001001001010;

			 118: data_out = 64'b1011111111011110000010111101001001110001111010010010100011100010;

			 119: data_out = 64'b1011111111011111000001110001111011101011101101010001000011111111;

			 120: data_out = 64'b1011111111011111111111111111111111111101110001100100110000000001;

			 121: data_out = 64'b1011111111100000011110110011000100011111111000011001010101111101;

			 122: data_out = 64'b1011111111100000111101010001100100111101100100010100011011000101;

			 123: data_out = 64'b1011111111100001011011011010111011010110010101011011011100000001;

			 124: data_out = 64'b1011111111100001111001001110100010000010111110000011011010100011;

			 125: data_out = 64'b1011111111100010010110101011110011110111011000111010000001100001;

			 126: data_out = 64'b1011111111100010110011110010001100000011010111011111001010001110;

			 127: data_out = 64'b1011111111100011010000100001000110010011001111111011110001100000;

			 128: data_out = 64'b1011111111100011101100110111111110110000101010010101000011000100;

			 129: data_out = 64'b1011111111100100001000110110010010000011001101011011000011001110;

			 130: data_out = 64'b1011111111100100100100011011011101010001001010110001111110001010;

			 131: data_out = 64'b1011111111100100111111100110111110000000001010010101000110100101;

			 132: data_out = 64'b1011111111100101011010011000010010010101110101010010101101000011;

			 133: data_out = 64'b1011111111100101110100101110111000111000100000011111111010000110;

			 134: data_out = 64'b1011111111100110001110101010010000101111110110000011110111011100;

			 135: data_out = 64'b1011111111100110101000001001111001100101011110011001010010101010;

			 136: data_out = 64'b1011111111100111000001001101010011100101101000100101100111011110;

			 137: data_out = 64'b1011111111100111011001110011111111011111110010000100111110111111;

			 138: data_out = 64'b1011111111100111110001111101011110100111001101101010010001111001;

			 139: data_out = 64'b1011111111101000001001101001010010110011101001110010011101011010;

			 140: data_out = 64'b1011111111101000100000110110111110100001110110001010011011000001;

			 141: data_out = 64'b1011111111101000110111100110000100110100001000100110101100010000;

			 142: data_out = 64'b1011111111101001001101110110001001010011000001001100001100011101;

			 143: data_out = 64'b1011111111101001100011100110110000001101101101101001011011000010;

			 144: data_out = 64'b1011111111101001111000110111011110011010101011111111010010101010;

			 145: data_out = 64'b1011111111101010001101100111111001011000001100011001000010000101;

			 146: data_out = 64'b1011111111101010100001110111100111001100110010010010011011110110;

			 147: data_out = 64'b1011111111101010110101100110001110100111110100101011110100000101;

			 148: data_out = 64'b1011111111101011001000110011010111000001111101101011000011101010;

			 149: data_out = 64'b1011111111101011011011011110101000011101101001001001001010000111;

			 150: data_out = 64'b1011111111101011101101100111101011100111100010101011100110111111;

			 151: data_out = 64'b1011111111101011111111001110001001110111000010101001000110000011;

			 152: data_out = 64'b1011111111101100010000010001101101001110101010011000111001111110;

			 153: data_out = 64'b1011111111101100100000110010000000011100011111101100100001111110;

			 154: data_out = 64'b1011111111101100110000101110101110111010100111010010111000100001;

			 155: data_out = 64'b1011111111101101000000000111100100101111011110100100101001111000;

			 156: data_out = 64'b1011111111101101001110111100001110101110010100011001010010010001;

			 157: data_out = 64'b1011111111101101011101001100011010010111100001000100000101000101;

			 158: data_out = 64'b1011111111101101101010110111110101111000111101011000111110110001;

			 159: data_out = 64'b1011111111101101110111111110010000001110011000111000100100111101;

			 160: data_out = 64'b1011111111101110000100011111011001000001101111000010111000111110;

			 161: data_out = 64'b1011111111101110010000011011000000101011011011110000100010001110;

			 162: data_out = 64'b1011111111101110011011110000111000010010101110110001110111000000;

			 163: data_out = 64'b1011111111101110100110100000110001101101111110010011101011011100;

			 164: data_out = 64'b1011111111101110110000101010011111100010111000101001001111010100;

			 165: data_out = 64'b1011111111101110111010001101110101000110110100111011000100110101;

			 166: data_out = 64'b1011111111101111000011001010100110011111000010111010011011011100;

			 167: data_out = 64'b1011111111101111001011100000101000100000111001111000111010110100;

			 168: data_out = 64'b1011111111101111010011001111110000110010000110100100001011111001;

			 169: data_out = 64'b1011111111101111011010010111110101101000111000000101001101111011;

			 170: data_out = 64'b1011111111101111100000111000101110001100001100000011001000000001;

			 171: data_out = 64'b1011111111101111100110110010010010010011111001101001000111100010;

			 172: data_out = 64'b1011111111101111101100000100011010101000111011101111011110000110;

			 173: data_out = 64'b1011111111101111110000101111000000100101011010000111010001111101;

			 174: data_out = 64'b1011111111101111110100110001111110010100110001101000110101101110;

			 175: data_out = 64'b1011111111101111111000001101001110110011111011100100011100111110;

			 176: data_out = 64'b1011111111101111111011000000101101110001010011110101100100110000;

			 177: data_out = 64'b1011111111101111111101001100010111101100111110011000001000000011;

			 178: data_out = 64'b1011111111101111111110110000001001111000101011011111111001101001;

			 179: data_out = 64'b1011111111101111111111101100000010010111111011010001111101110111;

			 180: data_out = 64'b1011111111110000000000000000000000000000000000000000000000000000;
			 
			 default: data_out = 64'd0;
		endcase
endmodule