module	SinDeg(input	signed	[7:0]		data_in,
					output	logic		[63:0]	data_out);

		always_comb
			case(data_in)
				-90: data_out = 64'b1011111111110000000000000000000000000000000000000000000000000000;

				-89: data_out = 64'b1011111111101111111111101100000010010111111100010110110110100000;

				-88: data_out = 64'b1011111111101111111110110000001001111000101101101001101001100101;

				-87: data_out = 64'b1011111111101111111101001100010111101101000001100110101100100110;

				-86: data_out = 64'b1011111111101111111011000000101101110001011000001000111001111001;

				-85: data_out = 64'b1011111111101111111000001101001110110100000000111100011101010100;

				-84: data_out = 64'b1011111111101111110100110001111110010100111000000101011010100100;

				-83: data_out = 64'b1011111111101111110000101111000000100101100001101000010011010001;

				-82: data_out = 64'b1011111111101111101100000100011010101001000100010100110010100000;

				-81: data_out = 64'b1011111111101111100110110010010010010100000011010010100100010100;

				-80: data_out = 64'b1011111111101111100000111000101110001100010110110000100001001001;

				-79: data_out = 64'b1011111111101111011010010111110101101001000011110110010110000011;

				-78: data_out = 64'b1011111111101111010011001111110000110010010011011000110100010100;

				-77: data_out = 64'b1011111111101111001011100000101000100001000111110000110011100010;

				-76: data_out = 64'b1011111111101111000011001010100110011111010001110101010011001001;

				-75: data_out = 64'b1011111111101110111010001101110101000111000100111000101000111011;

				-74: data_out = 64'b1011111111101110110000101010011111100011001001101001001011110111;

				-73: data_out = 64'b1011111111101110100110100000110001101110010000010101101011001111;

				-72: data_out = 64'b1011111111101110011011110000111000010011000001110101100011100011;

				-71: data_out = 64'b1011111111101110010000011011000000101011101111110101100011101111;

				-70: data_out = 64'b1011111111101110000100011111011001000010000100001000110110011011;

				-69: data_out = 64'b1011111111101101110111111110010000001110101110111111000100000000;

				-68: data_out = 64'b1011111111101101101010110111110101111001010100011111100011110110;

				-67: data_out = 64'b1011111111101101011101001100011010010111111001001010010011010110;

				-66: data_out = 64'b1011111111101101001110111100001110101110101101011110101011101100;

				-65: data_out = 64'b1011111111101101000000000111100100101111111000101000101111001001;

				-64: data_out = 64'b1011111111101100110000101110101110111011000010010101001001001000;

				-63: data_out = 64'b1011111111101100100000110010000000011100111011101100011100001010;

				-62: data_out = 64'b1011111111101100010000010001101101001111000111010101111010110100;

				-61: data_out = 64'b1011111111101011111111001110001001110111100000100010101001011100;

				-60: data_out = 64'b1011111111101011101101100111101011101000000001100001000111100110;

				-59: data_out = 64'b1011111111101011011011011110101000011110001000111010000001011110;

				-58: data_out = 64'b1011111111101011001000110011010111000010011110010110101010001001;

				-57: data_out = 64'b1011111111101010110101100110001110101000010110010001100000111010;

				-56: data_out = 64'b1011111111101010100001110111100111001101010100110001100101001001;

				-55: data_out = 64'b1011111111101010001101100111111001011000101111110000111100110010;

				-54: data_out = 64'b1011111111101001111000110111011110011011010000001111010010101001;

				-53: data_out = 64'b1011111111101001100011100110110000001110010010110000110011000100;

				-52: data_out = 64'b1011111111101001001101110110001001010011100111001010001110010000;

				-51: data_out = 64'b1011111111101000110111100110000100110100101111011010101000011010;

				-50: data_out = 64'b1011111111101000100000110110111110100010011101110011100001000100;

				-49: data_out = 64'b1011111111101000001001101001010010110100010010001111111011111101;

				-48: data_out = 64'b1011111111100111110001111101011110100111110110111011010110011110;

				-47: data_out = 64'b1011111111100111011001110011111111100000011100001000110110000100;

				-46: data_out = 64'b1011111111100111000001001101010011100110010011011011011100100101;

				-45: data_out = 64'b1011111111100110101000001001111001100110001010000000010000010110;

				-44: data_out = 64'b1011111111100110001110101010010000110000100010011011000111010110;

				-43: data_out = 64'b1011111111100101110100101110111000111001001101100110100100110100;

				-42: data_out = 64'b1011111111100101011010011000010010010110100011000111111010010000;

				-41: data_out = 64'b1011111111100100111111100110111110000000111000110111111101001100;

				-40: data_out = 64'b1011111111100100100100011011011101010001111010000001100100000011;

				-39: data_out = 64'b1011111111100100001000110110010010000011111101010110011101011110;

				-38: data_out = 64'b1011111111100011101100110111111110110001011010111011010101110110;

				-37: data_out = 64'b1011111111100011010000100001000110010100000001001100000000001100;

				-36: data_out = 64'b1011111111100010110011110010001100000100001001011000010111011010;

				-35: data_out = 64'b1011111111100010010110101011110011111000001011011011001110111010;

				-34: data_out = 64'b1011111111100001111001001110100010000011110001001011101001000111;

				-33: data_out = 64'b1011111111100001011011011010111011010111001001001001101011111101;

				-32: data_out = 64'b1011111111100000111101010001100100111110011000100111101011110111;

				-31: data_out = 64'b1011111111100000011110110011000100100000101101010000100110010100;

				-30: data_out = 64'b1011111111011111111111111111111111111111011100011001001100000000;

				-29: data_out = 64'b1011111111011111000001110001111011101101011001001001010110000100;

				-28: data_out = 64'b1011111111011110000010111101001001110011100111001100100101000000;

				-27: data_out = 64'b1011111111011101000011100010111000101010110000001111110010001000;

				-26: data_out = 64'b1011111111011100000011100100010111011010001111011110101010010110;

				-25: data_out = 64'b1011111111011011000011000010110101110110101110110110001011011101;

				-24: data_out = 64'b1011111111011010000001111111100100100000100011011110100101111100;

				-23: data_out = 64'b1011111111011001000000011011110100100010001001001110111111000000;

				-22: data_out = 64'b1011111111010111111110011000110111101110011101011100010000110101;

				-21: data_out = 64'b1011111111010110111011111000000000011111011000110101100110011101;

				-20: data_out = 64'b1011111111010101111000111010100001110100001000110000010011110100;

				-19: data_out = 64'b1011111111010100110101100001101111001111100111100101001001000010;

				-18: data_out = 64'b1011111111010011110001101110111100110110110100100001000010111111;

				-17: data_out = 64'b1011111111010010101101100011011111001111001010101011011010110100;

				-16: data_out = 64'b1011111111010001101001000000101011011100110111100011110111011000;

				-15: data_out = 64'b1011111111010000100100000111110111000001010000111001100100010101;

				-14: data_out = 64'b1011111111001110111101110100101111110010010011111100100110010001;

				-13: data_out = 64'b1011111111001100110010110011001000110110010000101110010110100100;

				-12: data_out = 64'b1011111111001010100111001101100110101011110000011010011110111111;

				-11: data_out = 64'b1011111111001000011011000110110111011100111111111111111100011010;

				-10: data_out = 64'b1011111111000110001110100001101001111101100111110111101001000010;

				-9: data_out = 64'b1011111111000100000001100000101101100111010001101101110110001010;

				-8: data_out = 64'b1011111111000001110100000110110010010110001101101100001001111000;

				-7: data_out = 64'b1011111110111111001100101101010001001011101101110000100011110100;

				-6: data_out = 64'b1011111110111010110000100110000010011010101110010111111010110100;

				-5: data_out = 64'b1011111110110110010011111101011010111000010101010100100000100000;

				-4: data_out = 64'b1011111110110001110110111000111101101101000100101101000110110011;

				-3: data_out = 64'b1011111110101010110010111100011101001000011011000110010111111100;

				-2: data_out = 64'b1011111110100001110111100101100011001001101000000011001110101110;

				-1: data_out = 64'b1011111110010001110111110000101100101011001100100010101001100011;

				0: data_out = 64'b0000000000000000000000000000000000000000000000000000000000000000;

				1: data_out = 64'b0011111110010001110111110000101100101011001100100010101001100011;

				2: data_out = 64'b0011111110100001110111100101100011001001101000000011001110101110;

				3: data_out = 64'b0011111110101010110010111100011101001000011011000110010111111100;

				4: data_out = 64'b0011111110110001110110111000111101101101000100101101000110110011;

				5: data_out = 64'b0011111110110110010011111101011010111000010101010100100000100000;

				6: data_out = 64'b0011111110111010110000100110000010011010101110010111111010110100;

				7: data_out = 64'b0011111110111111001100101101010001001011101101110000100011110100;

				8: data_out = 64'b0011111111000001110100000110110010010110001101101100001001111000;

				9: data_out = 64'b0011111111000100000001100000101101100111010001101101110110001010;

				10: data_out = 64'b0011111111000110001110100001101001111101100111110111101001000010;

				11: data_out = 64'b0011111111001000011011000110110111011100111111111111111100011010;

				12: data_out = 64'b0011111111001010100111001101100110101011110000011010011110111111;

				13: data_out = 64'b0011111111001100110010110011001000110110010000101110010110100100;

				14: data_out = 64'b0011111111001110111101110100101111110010010011111100100110010001;

				15: data_out = 64'b0011111111010000100100000111110111000001010000111001100100010101;

				16: data_out = 64'b0011111111010001101001000000101011011100110111100011110111011000;

				17: data_out = 64'b0011111111010010101101100011011111001111001010101011011010110100;

				18: data_out = 64'b0011111111010011110001101110111100110110110100100001000010111111;

				19: data_out = 64'b0011111111010100110101100001101111001111100111100101001001000010;

				20: data_out = 64'b0011111111010101111000111010100001110100001000110000010011110100;

				21: data_out = 64'b0011111111010110111011111000000000011111011000110101100110011101;

				22: data_out = 64'b0011111111010111111110011000110111101110011101011100010000110101;

				23: data_out = 64'b0011111111011001000000011011110100100010001001001110111111000000;

				24: data_out = 64'b0011111111011010000001111111100100100000100011011110100101111100;

				25: data_out = 64'b0011111111011011000011000010110101110110101110110110001011011101;

				26: data_out = 64'b0011111111011100000011100100010111011010001111011110101010010110;

				27: data_out = 64'b0011111111011101000011100010111000101010110000001111110010001000;

				28: data_out = 64'b0011111111011110000010111101001001110011100111001100100101000000;

				29: data_out = 64'b0011111111011111000001110001111011101101011001001001010110000100;

				30: data_out = 64'b0011111111011111111111111111111111111111011100011001001100000000;

				31: data_out = 64'b0011111111100000011110110011000100100000101101010000100110010100;

				32: data_out = 64'b0011111111100000111101010001100100111110011000100111101011110111;

				33: data_out = 64'b0011111111100001011011011010111011010111001001001001101011111101;

				34: data_out = 64'b0011111111100001111001001110100010000011110001001011101001000111;

				35: data_out = 64'b0011111111100010010110101011110011111000001011011011001110111010;

				36: data_out = 64'b0011111111100010110011110010001100000100001001011000010111011010;

				37: data_out = 64'b0011111111100011010000100001000110010100000001001100000000001100;

				38: data_out = 64'b0011111111100011101100110111111110110001011010111011010101110110;

				39: data_out = 64'b0011111111100100001000110110010010000011111101010110011101011110;

				40: data_out = 64'b0011111111100100100100011011011101010001111010000001100100000011;

				41: data_out = 64'b0011111111100100111111100110111110000000111000110111111101001100;

				42: data_out = 64'b0011111111100101011010011000010010010110100011000111111010010000;

				43: data_out = 64'b0011111111100101110100101110111000111001001101100110100100110100;

				44: data_out = 64'b0011111111100110001110101010010000110000100010011011000111010110;

				45: data_out = 64'b0011111111100110101000001001111001100110001010000000010000010110;

				46: data_out = 64'b0011111111100111000001001101010011100110010011011011011100100101;

				47: data_out = 64'b0011111111100111011001110011111111100000011100001000110110000100;

				48: data_out = 64'b0011111111100111110001111101011110100111110110111011010110011110;

				49: data_out = 64'b0011111111101000001001101001010010110100010010001111111011111101;

				50: data_out = 64'b0011111111101000100000110110111110100010011101110011100001000100;

				51: data_out = 64'b0011111111101000110111100110000100110100101111011010101000011010;

				52: data_out = 64'b0011111111101001001101110110001001010011100111001010001110010000;

				53: data_out = 64'b0011111111101001100011100110110000001110010010110000110011000100;

				54: data_out = 64'b0011111111101001111000110111011110011011010000001111010010101001;

				55: data_out = 64'b0011111111101010001101100111111001011000101111110000111100110010;

				56: data_out = 64'b0011111111101010100001110111100111001101010100110001100101001001;

				57: data_out = 64'b0011111111101010110101100110001110101000010110010001100000111010;

				58: data_out = 64'b0011111111101011001000110011010111000010011110010110101010001001;

				59: data_out = 64'b0011111111101011011011011110101000011110001000111010000001011110;

				60: data_out = 64'b0011111111101011101101100111101011101000000001100001000111100110;

				61: data_out = 64'b0011111111101011111111001110001001110111100000100010101001011100;

				62: data_out = 64'b0011111111101100010000010001101101001111000111010101111010110100;

				63: data_out = 64'b0011111111101100100000110010000000011100111011101100011100001010;

				64: data_out = 64'b0011111111101100110000101110101110111011000010010101001001001000;

				65: data_out = 64'b0011111111101101000000000111100100101111111000101000101111001001;

				66: data_out = 64'b0011111111101101001110111100001110101110101101011110101011101100;

				67: data_out = 64'b0011111111101101011101001100011010010111111001001010010011010110;

				68: data_out = 64'b0011111111101101101010110111110101111001010100011111100011110110;

				69: data_out = 64'b0011111111101101110111111110010000001110101110111111000100000000;

				70: data_out = 64'b0011111111101110000100011111011001000010000100001000110110011011;

				71: data_out = 64'b0011111111101110010000011011000000101011101111110101100011101111;

				72: data_out = 64'b0011111111101110011011110000111000010011000001110101100011100011;

				73: data_out = 64'b0011111111101110100110100000110001101110010000010101101011001111;

				74: data_out = 64'b0011111111101110110000101010011111100011001001101001001011110111;

				75: data_out = 64'b0011111111101110111010001101110101000111000100111000101000111011;

				76: data_out = 64'b0011111111101111000011001010100110011111010001110101010011001001;

				77: data_out = 64'b0011111111101111001011100000101000100001000111110000110011100010;

				78: data_out = 64'b0011111111101111010011001111110000110010010011011000110100010100;

				79: data_out = 64'b0011111111101111011010010111110101101001000011110110010110000011;

				80: data_out = 64'b0011111111101111100000111000101110001100010110110000100001001001;

				81: data_out = 64'b0011111111101111100110110010010010010100000011010010100100010100;

				82: data_out = 64'b0011111111101111101100000100011010101001000100010100110010100000;

				83: data_out = 64'b0011111111101111110000101111000000100101100001101000010011010001;

				84: data_out = 64'b0011111111101111110100110001111110010100111000000101011010100100;

				85: data_out = 64'b0011111111101111111000001101001110110100000000111100011101010100;

				86: data_out = 64'b0011111111101111111011000000101101110001011000001000111001111001;

				87: data_out = 64'b0011111111101111111101001100010111101101000001100110101100100110;

				88: data_out = 64'b0011111111101111111110110000001001111000101101101001101001100101;

				89: data_out = 64'b0011111111101111111111101100000010010111111100010110110110100000;

				90: data_out = 64'b0011111111110000000000000000000000000000000000000000000000000000;

		endcase
endmodule