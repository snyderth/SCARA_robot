
module Atan2 (
	areset,
	clk,
	q,
	x,
	y);	

	input		areset;
	input		clk;
	output	[12:0]	q;
	input	[31:0]	x;
	input	[31:0]	y;
endmodule
