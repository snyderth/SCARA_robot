module	CosDeg(input	signed	[7:0]		data_in,
					output	logic		[63:0]	data_out);

		always_comb
			case(data_in)
				-90: data_out = 64'b0011111000011110110101100000101000010001101001100010011000110011;

				-89: data_out = 64'b0011111110010001110111110000101101001010000001110000000001011000;

				-88: data_out = 64'b0011111110100001110111100101100011011001000010001101000011111101;

				-87: data_out = 64'b0011111110101010110010111100011101010111110100100000001000100101;

				-86: data_out = 64'b0011111110110001110110111000111101110100110000111000010101110110;

				-85: data_out = 64'b0011111110110110010011111101011011000000000000110100100000001100;

				-84: data_out = 64'b0011111110111010110000100110000010100010011001000011000110001001;

				-83: data_out = 64'b0011111110111111001100101101010001010011010111011101010110010111;

				-82: data_out = 64'b0011111111000001110100000110110010011010000001111110100101011000;

				-81: data_out = 64'b0011111111000100000001100000101101101011000101010111100010111110;

				-80: data_out = 64'b0011111111000110001110100001101010000001011010110011110111001010;

				-79: data_out = 64'b0011111111001000011011000110110111100000110010001001111100101111;

				-78: data_out = 64'b0011111111001010100111001101100110101111100001101101100011011000;

				-77: data_out = 64'b0011111111001100110010110011001000111010000001000101110010000110;

				-76: data_out = 64'b0011111111001110111101110100101111110110000011010011101100111001;

				-75: data_out = 64'b0011111111010000100100000111110111000011001000000010100111111000;

				-74: data_out = 64'b0011111111010001101001000000101011011110101110001000000110100000;

				-73: data_out = 64'b0011111111010010101101100011011111010001000000101000100001101000;

				-72: data_out = 64'b0011111111010011110001101110111100111000101001110100101110010010;

				-71: data_out = 64'b0011111111010100110101100001101111010001011100001101000110100001;

				-70: data_out = 64'b0011111111010101111000111010100001110101111100101010010001110110;

				-69: data_out = 64'b0011111111010110111011111000000000100001001011111111010100100010;

				-68: data_out = 64'b0011111111010111111110011000110111110000001111110011011111001101;

				-67: data_out = 64'b0011111111011001000000011011110100100011111010110001011111000110;

				-66: data_out = 64'b0011111111011010000001111111100100100010010100001010001001111010;

				-65: data_out = 64'b0011111111011011000011000010110101111000011110101000100110111000;

				-64: data_out = 64'b0011111111011100000011100100010111011011111110010101110001101011;

				-63: data_out = 64'b0011111111011101000011100010111000101100011110001001011011000110;

				-62: data_out = 64'b0011111111011110000010111101001001110101010100000110100110011011;

				-61: data_out = 64'b0011111111011111000001110001111011101111000101000001101000000101;

				-60: data_out = 64'b0011111111100000000000000000000000000000100011100110110100000000;

				-59: data_out = 64'b0011111111100000011110110011000100100001100010000111110110101100;

				-58: data_out = 64'b0011111111100000111101010001100100111111001100111010111100101000;

				-57: data_out = 64'b0011111111100001011011011010111011010111111100110111111011110111;

				-56: data_out = 64'b0011111111100001111001001110100010000100100100010011110111101001;

				-55: data_out = 64'b0011111111100010010110101011110011111000111101111100011100010010;

				-54: data_out = 64'b0011111111100010110011110010001100000100111011010001100100100100;

				-53: data_out = 64'b0011111111100011010000100001000110010100110010011100001110111000;

				-52: data_out = 64'b0011111111100011101100110111111110110010001011100001101000101000;

				-51: data_out = 64'b0011111111100100001000110110010010000100101101010001110111101101;

				-50: data_out = 64'b0011111111100100100100011011011101010010101001010001001001111101;

				-49: data_out = 64'b0011111111100100111111100110111110000001100111011010110011110010;

				-48: data_out = 64'b0011111111100101011010011000010010010111010000111101000111100000;

				-47: data_out = 64'b0011111111100101110100101110111000111001111010101101001111100000;

				-46: data_out = 64'b0011111111100110001110101010010000110001001110110010010111001110;

				-45: data_out = 64'b0011111111100110101000001001111001100110110101100111001110000100;

				-44: data_out = 64'b0011111111100111000001001101010011100110111110010001010001101100;

				-43: data_out = 64'b0011111111100111011001110011111111100001000110001100101101001010;

				-42: data_out = 64'b0011111111100111110001111101011110101000100000001100011011000010;

				-41: data_out = 64'b0011111111101000001001101001010010110100111010101101011010100001;

				-40: data_out = 64'b0011111111101000100000110110111110100011000101011100100111001010;

				-39: data_out = 64'b0011111111101000110111100110000100110101010110001110100100100011;

				-38: data_out = 64'b0011111111101001001101110110001001010100001101001000010000000001;

				-37: data_out = 64'b0011111111101001100011100110110000001110110111111000001011000101;

				-36: data_out = 64'b0011111111101001111000110111011110011011110100011111010010100111;

				-35: data_out = 64'b0011111111101010001101100111111001011001010011001000110111011111;

				-34: data_out = 64'b0011111111101010100001110111100111001101110111010000101110011100;

				-33: data_out = 64'b0011111111101010110101100110001110101000110111110111001101101111;

				-32: data_out = 64'b0011111111101011001000110011010111000010111111000010010000101000;

				-31: data_out = 64'b0011111111101011011011011110101000011110101000101010111000110110;

				-30: data_out = 64'b0011111111101011101101100111101011101000100000010110101000001101;

				-29: data_out = 64'b0011111111101011111111001110001001110111111110011100001100110100;

				-28: data_out = 64'b0011111111101100010000010001101101001111100100010010111011101011;

				-27: data_out = 64'b0011111111101100100000110010000000011101010111101100010110010111;

				-26: data_out = 64'b0011111111101100110000101110101110111011011101010111011001101110;

				-25: data_out = 64'b0011111111101101000000000111100100110000010010101100110100011010;

				-24: data_out = 64'b0011111111101101001110111100001110101111000110100100000101000111;

				-23: data_out = 64'b0011111111101101011101001100011010011000010001010000100001101001;

				-22: data_out = 64'b0011111111101101101010110111110101111001101011100110001000111011;

				-21: data_out = 64'b0011111111101101110111111110010000001111000101000101100011000100;

				-20: data_out = 64'b0011111111101110000100011111011001000010011001001110110011110111;

				-19: data_out = 64'b0011111111101110010000011011000000101100000011111010100101010001;

				-18: data_out = 64'b0011111111101110011011110000111000010011010100111001010000000110;

				-17: data_out = 64'b0011111111101110100110100000110001101110100010010111101011000010;

				-16: data_out = 64'b0011111111101110110000101010011111100011011010101001001000011010;

				-15: data_out = 64'b0011111111101110111010001101110101000111010100110110001101000000;

				-14: data_out = 64'b0011111111101111000011001010100110011111100000110000001010110110;

				-13: data_out = 64'b0011111111101111001011100000101000100001010101101000101100010000;

				-12: data_out = 64'b0011111111101111010011001111110000110010100000001101011100101110;

				-11: data_out = 64'b0011111111101111011010010111110101101001001111100111011110001010;

				-10: data_out = 64'b0011111111101111100000111000101110001100100001011101111010010001;

				-9: data_out = 64'b0011111111101111100110110010010010010100001100111100000001000111;

				-8: data_out = 64'b0011111111101111101100000100011010101001001100111010000110111010;

				-7: data_out = 64'b0011111111101111110000101111000000100101101001001001010100100110;

				-6: data_out = 64'b0011111111101111110100110001111110010100111110100001111111011011;

				-5: data_out = 64'b0011111111101111111000001101001110110100000110010100011101101010;

				-4: data_out = 64'b0011111111101111111011000000101101110001011100011100001111000001;

				-3: data_out = 64'b0011111111101111111101001100010111101101000100110101010001001001;

				-2: data_out = 64'b0011111111101111111110110000001001111000101111110011011001100001;

				-1: data_out = 64'b0011111111101111111111101100000010010111111101011011101111001001;

				0: data_out = 64'b0011111111110000000000000000000000000000000000000000000000000000;

				1: data_out = 64'b0011111111101111111111101100000010010111111101011011101111001001;

				2: data_out = 64'b0011111111101111111110110000001001111000101111110011011001100001;

				3: data_out = 64'b0011111111101111111101001100010111101101000100110101010001001001;

				4: data_out = 64'b0011111111101111111011000000101101110001011100011100001111000001;

				5: data_out = 64'b0011111111101111111000001101001110110100000110010100011101101010;

				6: data_out = 64'b0011111111101111110100110001111110010100111110100001111111011011;

				7: data_out = 64'b0011111111101111110000101111000000100101101001001001010100100110;

				8: data_out = 64'b0011111111101111101100000100011010101001001100111010000110111010;

				9: data_out = 64'b0011111111101111100110110010010010010100001100111100000001000111;

				10: data_out = 64'b0011111111101111100000111000101110001100100001011101111010010001;

				11: data_out = 64'b0011111111101111011010010111110101101001001111100111011110001010;

				12: data_out = 64'b0011111111101111010011001111110000110010100000001101011100101110;

				13: data_out = 64'b0011111111101111001011100000101000100001010101101000101100010000;

				14: data_out = 64'b0011111111101111000011001010100110011111100000110000001010110110;

				15: data_out = 64'b0011111111101110111010001101110101000111010100110110001101000000;

				16: data_out = 64'b0011111111101110110000101010011111100011011010101001001000011010;

				17: data_out = 64'b0011111111101110100110100000110001101110100010010111101011000010;

				18: data_out = 64'b0011111111101110011011110000111000010011010100111001010000000110;

				19: data_out = 64'b0011111111101110010000011011000000101100000011111010100101010001;

				20: data_out = 64'b0011111111101110000100011111011001000010011001001110110011110111;

				21: data_out = 64'b0011111111101101110111111110010000001111000101000101100011000100;

				22: data_out = 64'b0011111111101101101010110111110101111001101011100110001000111011;

				23: data_out = 64'b0011111111101101011101001100011010011000010001010000100001101001;

				24: data_out = 64'b0011111111101101001110111100001110101111000110100100000101000111;

				25: data_out = 64'b0011111111101101000000000111100100110000010010101100110100011010;

				26: data_out = 64'b0011111111101100110000101110101110111011011101010111011001101110;

				27: data_out = 64'b0011111111101100100000110010000000011101010111101100010110010111;

				28: data_out = 64'b0011111111101100010000010001101101001111100100010010111011101011;

				29: data_out = 64'b0011111111101011111111001110001001110111111110011100001100110100;

				30: data_out = 64'b0011111111101011101101100111101011101000100000010110101000001101;

				31: data_out = 64'b0011111111101011011011011110101000011110101000101010111000110110;

				32: data_out = 64'b0011111111101011001000110011010111000010111111000010010000101000;

				33: data_out = 64'b0011111111101010110101100110001110101000110111110111001101101111;

				34: data_out = 64'b0011111111101010100001110111100111001101110111010000101110011100;

				35: data_out = 64'b0011111111101010001101100111111001011001010011001000110111011111;

				36: data_out = 64'b0011111111101001111000110111011110011011110100011111010010100111;

				37: data_out = 64'b0011111111101001100011100110110000001110110111111000001011000101;

				38: data_out = 64'b0011111111101001001101110110001001010100001101001000010000000001;

				39: data_out = 64'b0011111111101000110111100110000100110101010110001110100100100011;

				40: data_out = 64'b0011111111101000100000110110111110100011000101011100100111001010;

				41: data_out = 64'b0011111111101000001001101001010010110100111010101101011010100001;

				42: data_out = 64'b0011111111100111110001111101011110101000100000001100011011000010;

				43: data_out = 64'b0011111111100111011001110011111111100001000110001100101101001010;

				44: data_out = 64'b0011111111100111000001001101010011100110111110010001010001101100;

				45: data_out = 64'b0011111111100110101000001001111001100110110101100111001110000100;

				46: data_out = 64'b0011111111100110001110101010010000110001001110110010010111001110;

				47: data_out = 64'b0011111111100101110100101110111000111001111010101101001111100000;

				48: data_out = 64'b0011111111100101011010011000010010010111010000111101000111100000;

				49: data_out = 64'b0011111111100100111111100110111110000001100111011010110011110010;

				50: data_out = 64'b0011111111100100100100011011011101010010101001010001001001111101;

				51: data_out = 64'b0011111111100100001000110110010010000100101101010001110111101101;

				52: data_out = 64'b0011111111100011101100110111111110110010001011100001101000101000;

				53: data_out = 64'b0011111111100011010000100001000110010100110010011100001110111000;

				54: data_out = 64'b0011111111100010110011110010001100000100111011010001100100100100;

				55: data_out = 64'b0011111111100010010110101011110011111000111101111100011100010010;

				56: data_out = 64'b0011111111100001111001001110100010000100100100010011110111101001;

				57: data_out = 64'b0011111111100001011011011010111011010111111100110111111011110111;

				58: data_out = 64'b0011111111100000111101010001100100111111001100111010111100101000;

				59: data_out = 64'b0011111111100000011110110011000100100001100010000111110110101100;

				60: data_out = 64'b0011111111100000000000000000000000000000100011100110110100000000;

				61: data_out = 64'b0011111111011111000001110001111011101111000101000001101000000101;

				62: data_out = 64'b0011111111011110000010111101001001110101010100000110100110011011;

				63: data_out = 64'b0011111111011101000011100010111000101100011110001001011011000110;

				64: data_out = 64'b0011111111011100000011100100010111011011111110010101110001101011;

				65: data_out = 64'b0011111111011011000011000010110101111000011110101000100110111000;

				66: data_out = 64'b0011111111011010000001111111100100100010010100001010001001111010;

				67: data_out = 64'b0011111111011001000000011011110100100011111010110001011111000110;

				68: data_out = 64'b0011111111010111111110011000110111110000001111110011011111001101;

				69: data_out = 64'b0011111111010110111011111000000000100001001011111111010100100010;

				70: data_out = 64'b0011111111010101111000111010100001110101111100101010010001110110;

				71: data_out = 64'b0011111111010100110101100001101111010001011100001101000110100001;

				72: data_out = 64'b0011111111010011110001101110111100111000101001110100101110010010;

				73: data_out = 64'b0011111111010010101101100011011111010001000000101000100001101000;

				74: data_out = 64'b0011111111010001101001000000101011011110101110001000000110100000;

				75: data_out = 64'b0011111111010000100100000111110111000011001000000010100111111000;

				76: data_out = 64'b0011111111001110111101110100101111110110000011010011101100111001;

				77: data_out = 64'b0011111111001100110010110011001000111010000001000101110010000110;

				78: data_out = 64'b0011111111001010100111001101100110101111100001101101100011011000;

				79: data_out = 64'b0011111111001000011011000110110111100000110010001001111100101111;

				80: data_out = 64'b0011111111000110001110100001101010000001011010110011110111001010;

				81: data_out = 64'b0011111111000100000001100000101101101011000101010111100010111110;

				82: data_out = 64'b0011111111000001110100000110110010011010000001111110100101011000;

				83: data_out = 64'b0011111110111111001100101101010001010011010111011101010110010111;

				84: data_out = 64'b0011111110111010110000100110000010100010011001000011000110001001;

				85: data_out = 64'b0011111110110110010011111101011011000000000000110100100000001100;

				86: data_out = 64'b0011111110110001110110111000111101110100110000111000010101110110;

				87: data_out = 64'b0011111110101010110010111100011101010111110100100000001000100101;

				88: data_out = 64'b0011111110100001110111100101100011011001000010001101000011111101;

				89: data_out = 64'b0011111110010001110111110000101101001010000001110000000001011000;

				90: data_out = 64'b0011111000011110110101100000101000010001101001100010011000110011;

		endcase
endmodule