// megafunction wizard: %ALTFP_SQRT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altfp_sqrt 

// ============================================================
// File Name: SqRoot.v
// Megafunction Name(s):
// 			altfp_sqrt
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 19.1.0 Build 670 09/22/2019 SJ Lite Edition
// ************************************************************


//Copyright (C) 2019  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and any partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details, at
//https://fpgasoftware.intel.com/eula.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module SqRoot (
	clk_en,
	clock,
	data,
	result);

	input	  clk_en;
	input	  clock;
	input	[63:0]  data;
	output	[63:0]  result;

	wire [63:0] sub_wire0;
	wire [63:0] result = sub_wire0[63:0];

	altfp_sqrt	altfp_sqrt_component (
				.clk_en (clk_en),
				.clock (clock),
				.data (data),
				.result (sub_wire0));
	defparam
		altfp_sqrt_component.pipeline = 30,
		altfp_sqrt_component.rounding = "TO_NEAREST",
		altfp_sqrt_component.width_exp = 11,
		altfp_sqrt_component.width_man = 52;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: FPM_FORMAT NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: PIPELINE NUMERIC "30"
// Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
// Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "11"
// Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "52"
// Retrieval info: USED_PORT: clk_en 0 0 0 0 INPUT NODEFVAL "clk_en"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: data 0 0 64 0 INPUT NODEFVAL "data[63..0]"
// Retrieval info: USED_PORT: result 0 0 64 0 OUTPUT NODEFVAL "result[63..0]"
// Retrieval info: CONNECT: @clk_en 0 0 0 0 clk_en 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 64 0 data 0 0 64 0
// Retrieval info: CONNECT: result 0 0 64 0 @result 0 0 64 0
// Retrieval info: GEN_FILE: TYPE_NORMAL SqRoot.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL SqRoot.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL SqRoot.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL SqRoot.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL SqRoot_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL SqRoot_bb.v FALSE
